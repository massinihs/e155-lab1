module (input logic reset_n, input logic [15:0] req, output logic [3:0] idx);

	always_comb begin
		casez(req)


		16'b0000 0000 0000 0001; idx = 4'b0001;
		16'b0000 0000 0000 0010; idx = 4'b0010;
		16'b0000 0000 0000 0100; idx = 4'b0011;
		16'b0000 0000 0000 1000; idx = 4'b0100;

		16'b0000 0000 0001 0000; idx = 4'b0101;
		16'b0000 0000 0010 0000; idx = 4'b0110;
		16'b0000 0000 0100 0000; idx = 4'b0111;
		16'b0000 0000 1000 0000; idx = 4'b1000;

		16'b0000 0001 0000 0000; idx = 4'b1001;
		16'b0000 0010 0000 0000; idx = 4'b1010;
		16'b0000 0100 0000 0000; idx = 4'b1011;
		16'b0000 1000 0000 0000; idx = 4'b1100;
		
		16'b0001 0000 0000 0000; idx = 4'b1101;
		16'b0010 0000 0000 0000; idx = 4'b1110;
		16'b0100 0000 0000 0000; idx = 4'b1111;


		endcase


	end



endmodule