//Massin Ihs
//mihs@g.hmc.edu
//9/8/2025
//Testbench to test the functionality of the 
//enable signals as well as the segment signals
 


`timescale 1ns/1ns
`default_nettype none
`define N_TV 8

module switcher_tb;

    // Inputs to DUT
    logic reset;
    logic [7:0] s;
    logic [6:0] seg;
    logic [1:0] enable;

    // Instantiate the DUT
   switcher dut (reset,s,seg,enable);
       

    initial begin
 

        reset = 1;
        s = 8'h2A; // A2

        #100;      // hold reset for 100 ns
        reset = 0;

        // change input after 2 ms
        #2000000;
        s = 8'h3C; // 3C


        #3000000;

        $finish;
    end



endmodule